//--------------------------------------------------------------------------------------------
// Module       : Interface
// Description  : Declaration of pin level signals as logic
//--------------------------------------------------------------------------------------------
interface spi_if;

  logic sclk;
  logic miso;
  logic mosi;
  logic ss;

endinterface
