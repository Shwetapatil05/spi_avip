//--------------------------------------------------------------------------------------------
// Module       : Slave Monitor BFM
// Description  : Connects the slave monitor bfm with the monitor proxy
//--------------------------------------------------------------------------------------------

module slave_monitor_bfm(spi_if intf);
  
  initial begin
    $display("Slave Monitor BFM");
  end

endmodule
